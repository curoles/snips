

//wire t = (select ? a : b);
`define MUX2(a, b) (select ? a : b)
