package helpers;

import stdtype::*;

//integer unsigned i = fill_with_1;
//
let fill_with_1() = '1;
let fill_with_0() = '0;
let fill_with_x() = 'x;
let fill_with_z() = 'z;

let get_parity(data) = ^data;

endpackage
