

module Bus ();

    parameter WIDTH = 1;

    wire [WIDTH-1:0] bus;

endmodule



